[aimspice]
[description]
1956
.include p18_cmos_models.inc
.include Photo-diode.inc

.param a=2

PhotoDiode_1 1 N1_1

*Vdd 1 0 1.8v
*Vex EXPOSE 0 1.8v
*Vnre NRE_R1 0 0v
*Ver ERASE 0 0v

*Ipd 1 N1_1 750p

*Photodiode 1*
*Mx DRAIN GATE SOURCE BULK*
M1_1 N1_1 EXPOSE N2_1 0 NMOS L=a*u W=a*2u
M2_1 N2_1 ERASE 0 0 NMOS L=a*u W=a*2u
M3_1 0 N2_1 N3_1 1 PMOS L=a*u W=a*2u
M4_1 N3_1 NRE_R1 OUT_1 1 PMOS L=a*u W=a*2u

CS_1 N2_1 0 3p


*Photodiode 2*
*Vnre NRE_R2 0 0v
*Ipd 1 N1_2 750p
*M1_2 N1_2 EXPOSE N2_2 0 NMOS L=a*u W=a*2u
*M2_2 N2_2 ERASE 0 0 NMOS L=a*u W=a*2u
*M3_2 0 N2_2 N3_2 1 PMOS L=a*u W=a*2u
*M4_2 N3_2 NRE_R2 OUT_2 1 PMOS L=a*u W=a*2u
*CS_2 N2_2 0 3p




.param Ipd_1 = 750p ! Photodiode current, range [50 pA, 750 pA]
.param VDD = 1.8 ! Supply voltage
.param EXPOSURETIME = 2m ! Exposure time, range [2 ms, 30 ms]

.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD = {EXPOSURETIME*10} ! Period for testbench sources
.param FS = 1k; ! Sampling clock frequency 
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_R1_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R1 signal
*.param NRE_R2_DLY = {4*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R2 signal
.param ERASE_DLY = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal

VDD 1 0 dc VDD
VEXPOSE EXPOSE 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE ERASE 0 dc 0 pulse(0 VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R1 NRE_R1 0 dc 0 pulse(VDD 0 NRE_R1_DLY TRF TRF CLK_PERIOD PERIOD)
*VNRE_R2 NRE_R2 0 dc 0  pulse(VDD 0 NRE_R2_DLY TRF TRF CLK_PERIOD PERIOD)

*.plot V(OUT1) V(OUT2) ! signals going to ADC
.plot V(OUT1) ! signals going to ADC

*.plot V(EXPOSE) V(NRE_R1) V(NRE_R2) V(ERASE)
.plot V(EXPOSE) V(NRE_R1)  V(ERASE)

.plot V(OUT_SAMPLED1)




[dc]
1
Vex
0
1.8
0.01
[tran]
0.001
0.06
X
X
0
[ana]
4 0
[end]
