
module Timer_counter(Initial, )