module basic_test_model();
    
    wire [0:3] pixels;

    initial begin
        

        $finish; // Done simulating
    end

endmodule